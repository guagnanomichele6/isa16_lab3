LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY ALU_CONTROL IS
	PORT (
		ALUop: IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		INSTR: IN STD_LOGIC_VECTOR(3 DOWNTO 0);	--func(6)&func3
		ALUctrl: OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
		);
END ENTITY;

ARCHITECTURE BEHAVIOR OF ALU_CONTROL IS

	SIGNAL AING: STD_LOGIC_VECTOR(5 DOWNTO 0);

BEGIN

	AING<=ALUop & INSTR;
	WITH AING SELECT ALUctrl <=
		"0010" WHEN "000000",--ADDI
		"0000" WHEN "000111",--ANDI
		"0011" WHEN "001101",--SRAI
		"0101" WHEN "010000",--U
		"0101" WHEN "010001",--U
		"0101" WHEN "010010",--U
		"0101" WHEN "010011",--U
		"0101" WHEN "010100",--U
		"0101" WHEN "010101",--U
		"0101" WHEN "010110",--U
		"0101" WHEN "010111",--U
		"0101" WHEN "011000",--U
		"0101" WHEN "011001",--U
		"0101" WHEN "011010",--U
		"0101" WHEN "011011",--U
		"0101" WHEN "011100",--U
		"0101" WHEN "011101",--U
		"0101" WHEN "011110",--U
		"0101" WHEN "011111",--U
		"0010" WHEN "100000",--ADD,ADDI,LW
		"0001" WHEN "100100",--XOR
		"0100" WHEN "100010",--SLT
		"1010" WHEN "110000",--J
		"1010" WHEN "110001",--J
		"1010" WHEN "110010",--J
		"1010" WHEN "110011",--J
		"1010" WHEN "110100",--J
		"1010" WHEN "110101",--J
		"1010" WHEN "110110",--J
		"1010" WHEN "110111",--J
		"1010" WHEN "111000",--J
		"1010" WHEN "111001",--J
		"1010" WHEN "111010",--J
		"1010" WHEN "111011",--J
		"1010" WHEN "111100",--J
		"1010" WHEN "111101",--J
		"1010" WHEN "111110",--J
		"1010" WHEN "111111",--J
		"0010" WHEN OTHERS;	--ADDI?(NOP)

END BEHAVIOR;
