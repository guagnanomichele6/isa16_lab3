library verilog;
use verilog.vl_types.all;
entity tb_riscv_abs is
end tb_riscv_abs;
