LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY WB IS
	PORT (	DM_READ_DATA_1:IN SIGNED(63 DOWNTO 0);
			ALU_RESULT_2: IN SIGNED(63 DOWNTO 0);
			MEMTOREG_3:IN STD_LOGIC;
			RF_WRITE_DATA: OUT SIGNED(63 DOWNTO 0)
		);
END WB;

ARCHITECTURE BEHAVIOR OF WB IS

BEGIN

WITH MEMTOREG_3 SELECT RF_WRITE_DATA<=
	DM_READ_DATA_1	WHEN '1',
	ALU_RESULT_2	WHEN OTHERS;

END BEHAVIOR;