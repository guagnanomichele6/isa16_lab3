LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY CU IS
	PORT (
		INSTRUCTION : IN STD_LOGIC_VECTOR(6 DOWNTO 0);
		CLK,RST,ZERO : IN STD_LOGIC;
		FUNC_1: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		RS1,RS2,RD2,RD3: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		FU_A,FU_B: OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
		ALU_OPERATION: OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		REG_WRITE_3, MEM_WRITE_2, MEM_READ_2,MEM_TO_REG_3,PC_SRC_3,ALU_SRC_1: OUT STD_LOGIC
	);
END CU;

ARCHITECTURE STRUCT OF CU IS

SIGNAL REG_WRITE,REG_WRITE_1,REG_WRITE_2,BRANCH_1,BRANCH_2,MEM_WRITE,MEM_WRITE_1:STD_LOGIC;
SIGNAL MEM_READ,MEM_READ_1,ZERO_1,MEM_TO_REG,MEM_TO_REG_1,MEM_TO_REG_2: STD_LOGIC;
SIGNAL ALU_SRC, BRANCH: STD_LOGIC;
SIGNAL ALU_OP,ALU_OP_1: STD_LOGIC_VECTOR(1 DOWNTO 0);
SIGNAL ALU_OUT: STD_LOGIC_VECTOR(7 DOWNTO 0);

COMPONENT FF IS
	PORT (
		D 				: IN STD_LOGIC;
		CLK,RST_N,EN 	: IN STD_LOGIC;
		Q				: OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT REG IS
	GENERIC (N:INTEGER);
	PORT (
		D 				: IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
		CLK,RST_N,EN 	: IN STD_LOGIC;
		Q				: OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0)
	);
END COMPONENT;

COMPONENT CONTROL IS
	PORT(
		INSTR: IN STD_LOGIC_VECTOR(6 DOWNTO 0);
		--BRANCH,MEM_READ,MEM_TO_REG,MEM_WRITE,ALU_SRC,REG_WRITE: OUT STD_LOGIC;
		--ALU_OP:  OUT STD_LOGIC_VECTOR(1 DOWNTO 0)
		ALU_OP: OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END COMPONENT;

COMPONENT ALU_CONTROL IS
	PORT(
		ALU_OP: IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		INSTR: IN STD_LOGIC_VECTOR(3 DOWNTO 0);--func(6)&func3
		ALU_OPERATION: OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END COMPONENT;

COMPONENT FORWARDING_UNIT IS
	PORT(
		RD_2, RD_3, RS_1, RS_2: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		FU_A, FU_B: OUT STD_LOGIC_VECTOR(1 DOWNTO 0)
	);
END COMPONENT;

BEGIN

--STAGE2
BRANCH<=ALU_OUT(7);
MEM_READ<=ALU_OUT(6);
MEM_TO_REG<=ALU_OUT(5);
ALU_OP<=ALU_OUT(4 DOWNTO 3);
MEM_WRITE<=ALU_OUT(2);
ALU_SRC<=ALU_OUT(1);
REG_WRITE<=ALU_OUT(0);
   CTRL: CONTROL
      PORT MAP (INSTRUCTION, ALU_OUT);


--REG ID/EX

   FF_MEMREAD: FF
      PORT MAP (MEM_READ,CLK,RST,'1',MEM_READ_1);

   FF_MEMWRITE: FF
      PORT MAP (MEM_WRITE,CLK,RST,'1',MEM_WRITE_1);

   FF_REGWRITE: FF
      PORT MAP (REG_WRITE,CLK,RST,'1',REG_WRITE_1);

   FF_BRANCH: FF
      PORT MAP (BRANCH,CLK,RST,'1',BRANCH_1);

   FF_MEMTOREG: FF
      PORT MAP (MEM_TO_REG,CLK,RST,'1',MEM_TO_REG_1);

   FF_ALUSRC: FF
      PORT MAP (ALU_SRC,CLK,RST,'1',ALU_SRC_1);

   REG_ALUOP: REG
      GENERIC MAP(2)
      PORT MAP (ALU_OP,CLK,RST,'1',ALU_OP_1);

--STAGE3

   FU: FORWARDING_UNIT
      PORT MAP (RD2,RD3,RS1,RS2,FU_A,FU_B);

   ALU_CTRL: ALU_CONTROL
      PORT MAP (ALU_OP_1,FUNC_1,ALU_OPERATION);

--REG EX/MEM

   FF_MEMREAD_1: FF
      PORT MAP (MEM_READ_1,CLK,RST,'1',MEM_READ_2);

   FF_MEMWRITE_1: FF
      PORT MAP (MEM_WRITE_1,CLK,RST,'1',MEM_WRITE_2);

   FF_BRANCH_1: FF
      PORT MAP (BRANCH_1,CLK,RST,'1',BRANCH_2);

   FF_MEMTOREG_1: FF
      PORT MAP (MEM_TO_REG_1,CLK,RST,'1',MEM_TO_REG_2);

   FF_REGWRITE_1: FF
      PORT MAP (REG_WRITE_1,CLK,RST,'1',REG_WRITE_2);

   FF_ZERO: FF
      PORT MAP (ZERO,CLK,RST,'1',ZERO_1);

--STAGE4

   PC_SRC_3<=BRANCH_2 AND ZERO_1;

--REG MEM/WB

   FF_REGWRITE_2: FF
      PORT MAP (REG_WRITE_2,CLK,RST,'1',REG_WRITE_3);

   FF_MEMTOREG_2: FF
      PORT MAP (MEM_TO_REG_2,CLK,RST,'1',MEM_TO_REG_3);

END STRUCT;