LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY COMPARATOR IS
	PORT(
		A, B: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		RES: OUT STD_LOGIC
	);
END ENTITY;

ARCHITECTURE BEHAVIOR OF COMPARATOR IS

SIGNAL ZERO: STD_LOGIC_VECTOR(4 DOWNTO 0);


BEGIN

	ZERO<= A XOR B;

WITH ZERO SELECT RES <=
    '1' WHEN "00000",
    '0' WHEN OTHERS;


END ARCHITECTURE;