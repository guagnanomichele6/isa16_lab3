LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY FULL_ADDER IS
	PORT (
		A 		: IN STD_LOGIC;
		B 		: IN STD_LOGIC;
		CIN		: IN STD_LOGIC;
		S 		: OUT STD_LOGIC;
		COUT 	: OUT STD_LOGIC
	);
END FULL_ADDER;

ARCHITECTURE STRUCT OF FULL_ADDER IS

BEGIN

	S 		<= A XOR B XOR CIN ;
	COUT 	<= (A AND B) OR (CIN AND A) OR (CIN AND B) ;

END STRUCT;