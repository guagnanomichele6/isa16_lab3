LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY DECODE IS
	PORT(	CLK,RST		 				: IN STD_LOGIC;
			PC_1						: IN UNSIGNED(63 DOWNTO 0);
			RD_3						: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
			INSTRUCTION_1 				: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
			RF_WRITE_DATA 				: IN SIGNED(63 DOWNTO 0);
			REGWRITE_3	  				: IN STD_LOGIC;
			FUNC						: OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
			RD							: OUT STD_LOGIC_vECTOR(4 DOWNTO 0);
			OPCODE						: OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
			PC_1_OUT					: OUT UNSIGNED(63 DOWNTO 0);
			IMM_OUT						: OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
			RF_READ_DATA1,RF_READ_DATA2 : OUT SIGNED(63 DOWNTO 0)
		);
END DECODE;

ARCHITECTURE BEHAVIOR OF DECODE IS

	COMPONENT REG_FILE IS
		PORT( 	WRITE_DATA 						: IN SIGNED (63 DOWNTO 0);
				REGWRITE,CLK,RST 				: IN STD_LOGIC;
				READ_REG1,READ_REG2,WRITE_REG 	: IN STD_LOGIC_VECTOR (4 DOWNTO 0); --32 regs
				READ_DATA1,READ_DATA2 			: OUT SIGNED (63 DOWNTO 0)
			);
	END COMPONENT;

	COMPONENT ImmGen IS	GENERIC (N : integer);
		PORT( 	A : IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
				B : OUT STD_LOGIC_VECTOR(2*N-1 DOWNTO 0)
			);
	END COMPONENT;

	SIGNAL READ_REG1,READ_REG2:STD_LOGIC_VECTOR(4 DOWNTO 0);

BEGIN

	OPCODE 		<= INSTRUCTION_1(6  DOWNTO 0);
	RD			<= INSTRUCTION_1(11 DOWNTO 7);
	READ_REG1 	<= INSTRUCTION_1(19 DOWNTO 15);
	READ_REG2 	<= INSTRUCTION_1(24 DOWNTO 20);
	FUNC		<= INSTRUCTION_1(30) & INSTRUCTION_1(14 DOWNTO 12);

	RF: REG_FILE
		PORT MAP (RF_WRITE_DATA,REGWRITE_3,CLK,RST,READ_REG1,READ_REG2,RD_3,RF_READ_DATA1,RF_READ_DATA2);

	IMM: IMMGEN
		GENERIC MAP(32)
		PORT MAP (INSTRUCTION_1,IMM_OUT);

	PC_1_OUT <= PC_1;

END ARCHITECTURE;