LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY CONTROL IS
	PORT(
		INSTR: IN STD_LOGIC_VECTOR(6 DOWNTO 0);
		--BRANCH,MEM_READ,MEM_TO_REG,MEM_WRITE,ALU_SRC,REG_WRITE: OUT STD_LOGIC;
		--ALU_OP:  OUT STD_LOGIC_VECTOR(1 DOWNTO 0)
		ALU_OP: OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END ENTITY;

ARCHITECTURE BEHAVIOR OF CONTROL IS

BEGIN

	--BRANCH<=INSTR(6);
	--MEM_READ<=INSTR(5);
	--MEM_TO_REG<=INSTR(4);
	WITH INSTR SELECT ALU_OP <=
	"01100111" WHEN "0000011", --LOAD --000 00 011
	"00000011" WHEN "0010011", --IMM --001 00 011
	"00000111" WHEN "0100011", --STORE
	"00010001" WHEN "0110011", --R  --000 10 001
	"10011000" WHEN "1100011", --BRANCH --100 11 000
	"00001011" WHEN "0110111", --U UPPER IMMEDIATE LUI  01
	"00001011" WHEN "0010111", --U UPPER IMMEDIATE AUIPC 01
	"00001011" WHEN "1101111", --J  
	"00000000" WHEN OTHERS; --00 is the op associated to I-type, I set others as NOP?

	--MEM_WRITE<=INSTR(2);
	--ALU_SRC<=INSTR(1);
	--REG_WRITE<=INSTR(0);

END ARCHITECTURE;