LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY ALU_CONTROL IS
	PORT(
		ALU_OP: IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		INSTR: IN STD_LOGIC_VECTOR(3 DOWNTO 0);--func(6)&func3
		ALU_OPERATION: OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END ENTITY;

ARCHITECTURE BEHAVIOR OF ALU_CONTROL IS

SIGNAL AING: STD_LOGIC_VECTOR(5 DOWNTO 0);
COMPONENT ADDER IS
        GENERIC(N:INTEGER);
	PORT (
		A 		: IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
		B 		: IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
		S 		: OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0);
		COUT 	: OUT STD_LOGIC
	);
END COMPONENT;

BEGIN

	AING<=ALU_OP&INSTR;
	WITH AING SELECT ALU_OPERATION <=
	"0010" WHEN "00----",--ADD
	"0110" WHEN "01----",--SUB
	"0010" WHEN "100000",--ADD
	"0110" WHEN "101000",--SUB
	"0000" WHEN "100111",--AND
	"0001" WHEN "100110", --OR
	"0111" WHEN "11----", --SUB, BRANCH
	"0010" WHEN OTHERS;--ADDI?(NOP)

END ARCHITECTURE;