LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY MUX_2TO1 IS
GENERIC (N:INTEGER);
    PORT ( SEL : IN  STD_LOGIC;
           A   : IN  STD_LOGIC_VECTOR (N-1 DOWNTO 0);
           B   : IN  STD_LOGIC_VECTOR (N-1 DOWNTO 0);
           X   : OUT STD_LOGIC_VECTOR (N-1 DOWNTO 0));
END MUX_2TO1;

ARCHITECTURE BEHAVIORAL OF MUX_2TO1 IS
BEGIN
    X <= A WHEN (SEL = '1') ELSE B;
END BEHAVIORAL;