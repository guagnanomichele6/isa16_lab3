LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY REG_FILE IS
	PORT(	WRITE_DATA 						: IN SIGNED (63 DOWNTO 0);
			REGWRITE, CLK, RST_N 			: IN STD_LOGIC;
			READ_REG1,READ_REG2,WRITE_REG 	: IN STD_LOGIC_VECTOR (4 DOWNTO 0); --32 regs
			READ_DATA1,READ_DATA2 			: OUT SIGNED (63 DOWNTO 0)
		);
END REG_FILE;

ARCHITECTURE BEHAVIOUR OF REG_FILE IS

	TYPE MEM_ARRAY IS ARRAY(0 TO 2**5-1) OF SIGNED (63 DOWNTO 0);
	SIGNAL MEM : MEM_ARRAY;

BEGIN

	PROCESS(CLK, RST_N)
		BEGIN
		IF (RST_N='0') THEN
			FOR i IN 0 TO 2**5-1 LOOP
				MEM(i)<=(OTHERS => '0');
			END LOOP;
		ELSIF (CLK'EVENT AND CLK='1' AND REGWRITE='1') THEN
			MEM(TO_INTEGER(UNSIGNED(WRITE_REG))) <= WRITE_DATA;
		END IF;
	END PROCESS;

	READ_DATA1 <= MEM(TO_INTEGER(UNSIGNED(READ_REG1)));
	READ_DATA2 <= MEM(TO_INTEGER(UNSIGNED(READ_REG2)));

END BEHAVIOUR;