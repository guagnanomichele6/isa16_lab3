LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY ADDER IS
GENERIC (N:INTEGER);
	PORT (
		A 		: IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
		B 		: IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
		CIN		: IN STD_LOGIC;
		S 		: OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0)
	);
END ADDER;

ARCHITECTURE STRUCT OF ADDER IS

SIGNAL COUT_SIGN: STD_LOGIC_VECTOR(N DOWNTO 0);

COMPONENT FULL_ADDER IS
	PORT (
		A 		: IN STD_LOGIC;
		B 		: IN STD_LOGIC;
		CIN		: IN STD_LOGIC;
		S 		: OUT STD_LOGIC;
		COUT 	: OUT STD_LOGIC
	);
END COMPONENT;

BEGIN
COUT_SIGN(0)<='0';
GEN_FA : FOR I IN 0 TO N-1 GENERATE 
   FA: FULL_ADDER PORT MAP(A(I),B(I),COUT_SIGN(I),S(I),COUT_SIGN(I+1));
END GENERATE GEN_FA;

END STRUCT;