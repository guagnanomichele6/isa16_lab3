LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY MEM IS 
					PORT(	ALU_RESULT_1:IN SIGNED(63 DOWNTO 0);
							DM_ADDRESS :OUT SIGNED(63 DOWNTO 0);
							RF_READ_DATA2_2: IN SIGNED(63 DOWNTO 0);
							DM_WRITE_DATA:OUT SIGNED(63 DOWNTO 0);
							DM_READ_DATA:IN SIGNED(63 DOWNTO 0);
							DM_READ_DATA_OUT: OUT SIGNED(63 DOWNTO 0);
							RD_2:IN STD_LOGIC_VECTOR(4 DOWNTO 0);
							RD_2_OUT:OUT STD_LOGIC_VECTOR(4 DOWNTO 0)
							 );	
END MEM;

ARCHITECTURE STRUCT OF MEM IS 

--DATA MEMORY IS IN THE TESTBENCH

BEGIN

DM_ADDRESS<=ALU_RESULT_1;
DM_WRITE_DATA<=RF_READ_DATA2_2;
DM_READ_DATA_OUT<=DM_READ_DATA;
RD_2_OUT<=RD_2;

END STRUCT;
