LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY RISCV_pipeline_abs IS
	PORT (
		CLK,RST_N: IN STD_LOGIC;
		INSTRUCTION: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		DM_READ_DATA: IN SIGNED(63 DOWNTO 0);
		IM_ADDRESS: OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
		MEMWRITE_OUT,MEMREAD_OUT: OUT STD_LOGIC;
		DM_ADDRESS: OUT SIGNED(63 DOWNTO 0);
		DM_WRITE_DATA: OUT SIGNED(63 DOWNTO 0)
		);
END ENTITY;

ARCHITECTURE STRUCT OF RISCV_pipeline_abs IS

	COMPONENT FETCH IS
		PORT (
			CLK,RST_N: IN STD_LOGIC;
			BRANCH_SUM:IN SIGNED(63 DOWNTO 0);
			PCsrc  : IN STD_LOGIC;
			PC_OUT : OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
			INSTRUCTION: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
			INSTRUCTION_OUT: OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
			);
	END COMPONENT;

	COMPONENT DECODE IS
		PORT (
			CLK,RST_N		 : IN STD_LOGIC;
			PC_1			 : IN UNSIGNED(63 DOWNTO 0);
			RD_3			 : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
			INSTRUCTION_1: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
			RF_WRITE_DATA: IN SIGNED(63 DOWNTO 0);
			REGWRITE_3	 : IN STD_LOGIC;
			FUNC			 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
			RD				 : OUT STD_LOGIC_vECTOR(4 DOWNTO 0);
			OPCODE		 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
			PC_1_OUT		 : OUT UNSIGNED(63 DOWNTO 0);
			IMM_OUT		 : OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
			RF_READ_DATA1,RF_READ_DATA2: OUT SIGNED(63 DOWNTO 0)
			);
	END COMPONENT;

	COMPONENT EXECUTE_abs IS
		PORT (
			PC_2,IMM_OUT_1:IN SIGNED(63 DOWNTO 0);
			RD_1: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
			READ_DATA1_1,READ_DATA2_1:IN SIGNED(63 DOWNTO 0);
			ALUctrl: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			ALUsrc1_1: IN STD_LOGIC;
			ALUsrc2_1: IN STD_LOGIC;
			ZERO: OUT STD_LOGIC;
			RD_1_OUT: OUT STD_LOGIC_VECTOR(4 DOWNTO 0);
			BRANCH_SUM: OUT SIGNED (63 DOWNTO 0);
			ALU_RESULT: OUT SIGNED(63 DOWNTO 0);
			RF_READ_DATA2_1_OUT: OUT SIGNED(63 DOWNTO 0)
			);
	END COMPONENT;

	COMPONENT MEM IS
		PORT (
			ALU_RESULT_1:IN SIGNED(63 DOWNTO 0);
			DM_ADDRESS :OUT SIGNED(63 DOWNTO 0);
			RF_READ_DATA2_2: IN SIGNED(63 DOWNTO 0);
			DM_WRITE_DATA:OUT SIGNED(63 DOWNTO 0);
			DM_READ_DATA:IN SIGNED(63 DOWNTO 0);
			DM_READ_DATA_OUT: OUT SIGNED(63 DOWNTO 0);
			RD_2:IN STD_LOGIC_VECTOR(4 DOWNTO 0);
			RD_2_OUT:OUT STD_LOGIC_VECTOR(4 DOWNTO 0)
			);
	END COMPONENT;

	COMPONENT WB IS
		PORT (
			DM_READ_DATA_1:IN SIGNED(63 DOWNTO 0);
			ALU_RESULT_2: IN SIGNED(63 DOWNTO 0);
			MEMTOREG_3:IN STD_LOGIC;
			RF_WRITE_DATA: OUT SIGNED(63 DOWNTO 0)
			);
	END COMPONENT;

	COMPONENT CONTROL IS
		PORT (
			OPCODE   : IN  STD_LOGIC_VECTOR(6 DOWNTO 0);
			BRANCH   : OUT STD_LOGIC;
			MEMREAD  : OUT STD_LOGIC;
			MEMTOREG : OUT STD_LOGIC;
			ALUop	   : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
			MEMWRITE : OUT STD_LOGIC;
			ALUsrc1  : OUT STD_LOGIC;
			ALUsrc2  : OUT STD_LOGIC;
			REGWRITE : OUT STD_LOGIC
			);
	END COMPONENT;

	COMPONENT ALU_CONTROL_abs IS
		PORT (
			ALUop: IN STD_LOGIC_VECTOR(1 DOWNTO 0);
			INSTR: IN STD_LOGIC_VECTOR(3 DOWNTO 0);	--func(6)&func3
			ALUctrl: OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
			);
	END COMPONENT;

	SIGNAL PCsrc															: STD_LOGIC;
	SIGNAL INSTRUCTION_OUT													: STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL INSTRUCTION_1													: STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL PC_OUT															: STD_LOGIC_VECTOR(63 DOWNTO 0);
	SIGNAL PC_1,PC_1_OUT													: UNSIGNED(63 DOWNTO 0);
	SIGNAL PC_2																: SIGNED(63 DOWNTO 0);
	SIGNAL FUNC,FUNC_1														: STD_LOGIC_VECTOR(3 DOWNTO 0);
	SIGNAL RD,RD_1,RD_1_OUT,RD_2,RD_2_OUT,RD_3								: STD_LOGIC_VECTOR(4 DOWNTO 0);
	SIGNAL RF_READ_DATA1,RF_READ_DATA1_1									: SIGNED (63 DOWNTO 0);
	SIGNAL RF_READ_DATA2,RF_READ_DATA2_1,RF_READ_DATA2_1_OUT,RF_READ_DATA2_2: SIGNED (63 DOWNTO 0);
	SIGNAL OPCODE															: STD_LOGIC_VECTOR(6 DOWNTO 0);
	SIGNAL IMM_OUT															: STD_LOGIC_VECTOR(63 DOWNTO 0);	-----------NON DEVE ESSERE SIGNED?
	SIGNAL IMM_OUT_1														: SIGNED(63 DOWNTO 0);
	SIGNAL REGWRITE,REGWRITE_1,REGWRITE_2,REGWRITE_3						: STD_LOGIC;
	SIGNAL ALUop,ALUop_1													: STD_LOGIC_VECTOR(1 DOWNTO 0);
	SIGNAL ALUsrc1,ALUsrc1_1												: STD_LOGIC;
	SIGNAL ALUsrc2,ALUsrc2_1												: STD_LOGIC;
	SIGNAL MEMTOREG,MEMTOREG_1,MEMTOREG_2,MEMTOREG_3						: STD_LOGIC;
	SIGNAL BRANCH,BRANCH_1,BRANCH_2											: STD_LOGIC;
	SIGNAL MEMREAD,MEMREAD_1,MEMREAD_2										: STD_LOGIC;
	SIGNAL MEMWRITE,MEMWRITE_1,MEMWRITE_2									: STD_LOGIC;
	SIGNAL ALUctrl															: STD_LOGIC_VECTOR(3 DOWNTO 0);
	SIGNAL ZERO,ZERO_1														: STD_LOGIC;
	SIGNAL BRANCH_SUM,BRANCH_SUM_1											: SIGNED(63 DOWNTO 0);
	SIGNAL ALU_RESULT,ALU_RESULT_1,ALU_RESULT_2								: SIGNED(63 DOWNTO 0);
	SIGNAL DM_READ_DATA_OUT,DM_READ_DATA_1,DM_WRITE_DATA_OUT				: SIGNED(63 DOWNTO 0);
	SIGNAL RF_WRITE_DATA													: SIGNED(63 DOWNTO 0);

BEGIN
	IM_ADDRESS		<= PC_OUT;
	MEMWRITE_OUT	<= MEMWRITE_2;
	MEMREAD_OUT		<= MEMREAD_2;

	IF_STAGE: FETCH
		PORT MAP (CLK,RST_N,BRANCH_SUM_1,PCsrc,PC_OUT,INSTRUCTION,INSTRUCTION_OUT);
	-------------------------------------------------------------------------------------------------------
	-- PIPELINE REGISTER stage 1
	PROCESS(CLK,RST_N)
	BEGIN
		IF (RST_N='0') THEN
			PC_1			<= (OTHERS=>'0');
			INSTRUCTION_1	<= (OTHERS=>'0');
		ELSIF (CLK'EVENT AND CLK='1') THEN
			PC_1			<= UNSIGNED(PC_OUT);
			INSTRUCTION_1	<= INSTRUCTION_OUT;
		END IF;
	END PROCESS;
	-------------------------------------------------------------------------------------------------------
	ID_STAGE: DECODE
		PORT MAP (CLK,RST_N,PC_1,RD_3,INSTRUCTION_1,RF_WRITE_DATA,REGWRITE_3,FUNC,RD,OPCODE,PC_1_OUT,IMM_OUT,RF_READ_DATA1,RF_READ_DATA2);
	ID_CTRL: CONTROL
		PORT MAP (OPCODE,BRANCH,MEMREAD,MEMTOREG,ALUop,MEMWRITE,ALUsrc1,ALUsrc2,REGWRITE);
	-------------------------------------------------------------------------------------------------------
	-- PIPELINE REGISTER stage 2
	PROCESS(CLK,RST_N)
	BEGIN
		IF (RST_N='0') THEN
			PC_2			<= (OTHERS=>'0');
			IMM_OUT_1		<= (OTHERS=>'0');
			FUNC_1			<= (OTHERS=>'0');
			RD_1			<= (OTHERS=>'0');
			RF_READ_DATA1_1	<= (OTHERS=>'0');
			RF_READ_DATA2_1	<= (OTHERS=>'0');

			BRANCH_1		<= '0';
			MEMREAD_1		<= '0';
			MEMTOREG_1		<= '0';
			ALUop_1			<= (OTHERS=>'0');
			MEMWRITE_1		<= '0';
			ALUsrc1_1		<= '0';
			ALUsrc2_1		<= '0';
			REGWRITE_1		<= '0';
		ELSIF (CLK'EVENT AND CLK='1') THEN
			PC_2			<= SIGNED(PC_1_OUT);
			IMM_OUT_1		<= SIGNED(IMM_OUT);
			FUNC_1			<= FUNC;
			RD_1			<= RD;
			RF_READ_DATA1_1	<= RF_READ_DATA1;
			RF_READ_DATA2_1	<= RF_READ_DATA2;

			BRANCH_1		<= BRANCH;
			MEMREAD_1		<= MEMREAD;
			MEMTOREG_1		<= MEMTOREG;
			ALUop_1			<= ALUop;
			MEMWRITE_1		<= MEMWRITE;
			ALUsrc1_1		<= ALUsrc1;
			ALUsrc2_1		<= ALUsrc2;
			REGWRITE_1		<= REGWRITE;
		END IF;
	END PROCESS;
	-------------------------------------------------------------------------------------------------------
	EX_STAGE: EXECUTE_abs
		PORT MAP (PC_2,IMM_OUT_1,RD_1,RF_READ_DATA1_1,RF_READ_DATA2_1,ALUctrl,ALUsrc1_1,ALUsrc2_1,ZERO,RD_1_OUT,BRANCH_SUM,ALU_RESULT,RF_READ_DATA2_1_OUT);
	EX_CTRL: ALU_CONTROL_abs
		PORT MAP (ALUop_1,FUNC_1,ALUctrl);
	-------------------------------------------------------------------------------------------------------
	--PIPELINE REGISTER stage 3
	PROCESS(CLK,RST_N)
	BEGIN
		IF (RST_N='0') THEN
			ALU_RESULT_1	<= (OTHERS=>'0');
			RF_READ_DATA2_2	<= (OTHERS=>'0');
			RD_2			<= (OTHERS=>'0');
			ZERO_1			<= '0';

			BRANCH_2		<= '0';
			MEMREAD_2		<= '0';
			MEMTOREG_2		<= '0';
			MEMWRITE_2		<= '0';
			REGWRITE_2		<= '0';
			BRANCH_SUM_1	<= (OTHERS=>'0');
		ELSIF (CLK'EVENT AND CLK='1') THEN
			ALU_RESULT_1	<= ALU_RESULT;
			RF_READ_DATA2_2	<= RF_READ_DATA2_1_OUT;
			RD_2			<= RD_1_OUT;
			ZERO_1			<= ZERO;

			BRANCH_2		<= BRANCH_1;
			MEMREAD_2		<= MEMREAD_1;
			MEMTOREG_2		<= MEMTOREG_1;
			MEMWRITE_2		<= MEMWRITE_1;
			REGWRITE_2		<= REGWRITE_1;
			BRANCH_SUM_1	<= BRANCH_SUM;
		END IF;
	END PROCESS;
	-------------------------------------------------------------------------------------------------------
	MEM_STAGE: MEM
		PORT MAP(ALU_RESULT_1,DM_ADDRESS,RF_READ_DATA2_2,DM_WRITE_DATA,DM_READ_DATA,DM_READ_DATA_OUT,RD_2,RD_2_OUT);
	PCsrc <= BRANCH_2 AND ZERO_1;
	-------------------------------------------------------------------------------------------------------
	--PIPELINE REGISTER stage 4
	PROCESS(CLK,RST_N)
	BEGIN
		IF (RST_N='0') THEN
			ALU_RESULT_2	<= (OTHERS=>'0');
			DM_READ_DATA_1	<= (OTHERS=>'0');
			RD_3			<= (OTHERS=>'0');

			MEMTOREG_3		<= '0';
			REGWRITE_3		<= '0';
		ELSIF (CLK'EVENT AND CLK='1') THEN
			ALU_RESULT_2	<= ALU_RESULT_1;
			DM_READ_DATA_1	<= DM_READ_DATA_OUT;
			RD_3			<= RD_2_OUT;

			MEMTOREG_3		<= MEMTOREG_2;
			REGWRITE_3		<= REGWRITE_2;
		END IF;
	END PROCESS;
	-------------------------------------------------------------------------------------------------------
	WB_STAGE: WB
		PORT MAP(DM_READ_DATA_1,ALU_RESULT_2,MEMTOREG_3,RF_WRITE_DATA);

END STRUCT;
