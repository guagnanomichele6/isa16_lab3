LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY DATAPATH IS
	PORT(
		CLK, RST, MUX_PC_SEL, MUX_ALU_SEL, MUX_WB_SEL, REGWRITE: IN STD_LOGIC;
		READ_DATA: IN SIGNED(63 DOWNTO 0);
		INSTR: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		ALU_OPERATION: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		RD2,RD3,RS1,RS2: OUT STD_LOGIC_VECTOR(4 DOWNTO 0);
		FU_A, FU_B: IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		ZERO: OUT STD_LOGIC;
		ALU_RESULT_1: OUT SIGNED(63 DOWNTO 0);
		READ_DATA1_3: OUT SIGNED(63 DOWNTO 0);
		OPCODE: OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
		FUNC_1: OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		PC_O: OUT STD_LOGIC_VECTOR(63 DOWNTO 0)
	);
END ENTITY;

ARCHITECTURE BEHAVIOR OF DATAPATH IS

SIGNAL SUM,SUM_1: STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL IMM_OUT,IMM_OUT1: STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL READ_DATA1,READ_DATA2,READ_DATA1_1,READ_DATA2_1,READ_DATA1_2, ALU_RESULT, ALU_RESULT_2,ALU_RESULT_1_SIGNAL: SIGNED(63 DOWNTO 0);
SIGNAL IMM_OUT1_SHIFTED: STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL MUX_WB_OUT,MUX_ALU_OUT,MUX_ALU_OUT_1,READ_DATA_1: SIGNED(63 DOWNTO 0);
SIGNAL PC,PC_SIGNAL,MUX_PC_OUT,PC_1,PC_2,PC_PLUS_4: STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL RD,RD_1,RD_2,RD_3,READ_REG1,READ_REG2,READ_REG1_1,READ_REG2_1: STD_LOGIC_VECTOR(4 DOWNTO 0);
SIGNAL FUNC: STD_LOGIC_VECTOR( 3 DOWNTO 0);
SIGNAL INSTRUCTION: STD_LOGIC_VECTOR(31 DOWNTO 0);


COMPONENT MUX_2TO1 IS
GENERIC (N:INTEGER);
    PORT ( SEL : IN  STD_LOGIC;
           A   : IN  STD_LOGIC_VECTOR (N-1 DOWNTO 0);
           B   : IN  STD_LOGIC_VECTOR (N-1 DOWNTO 0);
           X   : OUT STD_LOGIC_VECTOR (N-1 DOWNTO 0));
END COMPONENT;

COMPONENT MUX_3 IS
GENERIC (N:INTEGER);
    PORT ( SEL : IN  STD_LOGIC_VECTOR(1 DOWNTO 0);
           A   : IN  SIGNED (N-1 DOWNTO 0);
           B   : IN  SIGNED (N-1 DOWNTO 0);
           C   : IN  SIGNED (N-1 DOWNTO 0);
           X   : OUT SIGNED (N-1 DOWNTO 0));
END COMPONENT;

COMPONENT MUX_DATA IS
GENERIC (N:INTEGER);
    PORT ( SEL : IN  STD_LOGIC;
           A   : IN  SIGNED (N-1 DOWNTO 0);
           B   : IN  SIGNED (N-1 DOWNTO 0);
           X   : OUT SIGNED (N-1 DOWNTO 0));
END COMPONENT;

COMPONENT ImmGen IS
  GENERIC (N : integer);
 PORT (
		A : IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
		B : OUT STD_LOGIC_VECTOR(2*N-1 DOWNTO 0)
	);
END COMPONENT;

COMPONENT REG_FILE IS     
 PORT( WRITE_DATA : IN SIGNED (63 DOWNTO 0);
		 REGWRITE,CLK,RST : IN STD_LOGIC;
		 READ_REG1,READ_REG2,WRITE_REG : IN STD_LOGIC_VECTOR (4 DOWNTO 0); --32 regs
		 READ_DATA1,READ_DATA2 : OUT SIGNED (63 DOWNTO 0));
END COMPONENT;

COMPONENT ADDER IS
        GENERIC(N:INTEGER);
	PORT (
		A 		: IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
		B 		: IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
		CIN		: IN STD_LOGIC;
		S 		: OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0)
	);
END COMPONENT;

COMPONENT REG IS
	GENERIC (N:INTEGER);
	PORT (
		D 				: IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
		CLK,RST_N,EN 	: IN STD_LOGIC;
		Q				: OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0)
	);
END COMPONENT;

COMPONENT PC_REG IS
	PORT (
		D 				: IN STD_LOGIC_VECTOR(63 DOWNTO 0);
		CLK,RST_N,EN 	: IN STD_LOGIC;
		Q				: OUT STD_LOGIC_VECTOR(63 DOWNTO 0)
	);
END COMPONENT;

COMPONENT REG_DATA IS
	GENERIC (N:INTEGER);
	PORT (
		D 				: IN SIGNED(N-1 DOWNTO 0);
		CLK,RST_N,EN 	: IN STD_LOGIC;
		Q				: OUT SIGNED(N-1 DOWNTO 0)
	);
END COMPONENT;

COMPONENT ALU IS
	PORT(
		A: IN SIGNED(63 DOWNTO 0);
		B: IN SIGNED(63 DOWNTO 0);
		ALU_OPERATION: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		CLK				: IN STD_LOGIC;
		ZERO: OUT STD_LOGIC;
		ALU_RESULT: OUT SIGNED(63 DOWNTO 0)
	);
END COMPONENT;

COMPONENT SHIFT_REG_1 IS
  GENERIC (N : integer);
 PORT (
		D 				: IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
		CLK,RST_N,EN 	: IN STD_LOGIC;
		Q				: OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0)
	);
END COMPONENT;

BEGIN

--STAGE1
   MUX_PC: MUX_2TO1
      GENERIC MAP(64)
      PORT MAP (MUX_PC_SEL, SUM_1, PC_PLUS_4 ,MUX_PC_OUT);

   PREG_PC: REG
      GENERIC MAP(64)
      PORT MAP (MUX_PC_OUT,CLK,RST,'1',PC_SIGNAL);

   PC_ADD:  ADDER
      GENERIC MAP(64)
      PORT MAP(PC_SIGNAL,std_logic_vector(to_unsigned(4, 64)),'0',PC_PLUS_4);

--REG IF/ID
   PC<=PC_SIGNAL;
   PC_O<=PC;--(7 DOWNTO 0);

   REG_PC_IF: REG
      GENERIC MAP(64)
      PORT MAP (PC_SIGNAL,CLK,RST,'1',PC_1);

   REG_INSTR_IF: REG
      GENERIC MAP(32)
      PORT MAP (INSTR,CLK,RST,'1',INSTRUCTION);

--STAGE2

READ_REG1<=INSTRUCTION(19 DOWNTO 15);
READ_REG2<=INSTRUCTION(24 DOWNTO 20);
   RF: REG_FILE
      PORT MAP (MUX_WB_OUT,REGWRITE,CLK,RST,READ_REG1,READ_REG2,RD_3,READ_DATA1,READ_DATA2);   

   IMM: IMMGEN
      GENERIC MAP(32)
      PORT MAP (INSTRUCTION,IMM_OUT);

   OPCODE <= INSTRUCTION(6 DOWNTO 0);

   RD<=INSTRUCTION(11 DOWNTO 7);

--REG ID/EX

   REG_PC_ID: REG
      GENERIC MAP(64)
      PORT MAP (PC_1,CLK,RST,'1',PC_2);

   REG_READ_DATA1_ID: REG_DATA
      GENERIC MAP(64)
      PORT MAP (READ_DATA1,CLK,RST,'1',READ_DATA1_1);

   REG_READ_DATA2_ID: REG_DATA
      GENERIC MAP(64)
      PORT MAP (READ_DATA2,CLK,RST,'1',READ_DATA2_1);

   REG_IMMGEN_ID: REG
      GENERIC MAP(64)
      PORT MAP (IMM_OUT,CLK,RST,'1',IMM_OUT1);

   REG_READREAG1_ID: REG
      GENERIC MAP(5)
      PORT MAP (READ_REG1,CLK,RST,'1',READ_REG1_1);

   REG_READREAG2_ID: REG
      GENERIC MAP(5)
      PORT MAP (READ_REG2,CLK,RST,'1',READ_REG2_1);

   REG_RD_ID: REG
      GENERIC MAP(5)
      PORT MAP (RD,CLK,RST,'1',RD_1);

FUNC<=INSTR(30)&INSTR(14 DOWNTO 12);

   REG_FUNC_ID: REG
      GENERIC MAP(4)
      PORT MAP (FUNC,CLK,RST,'1',FUNC_1);

--STAGE3

   RD2<=RD_2;
   RD3<=RD_3;
   RS1<=READ_REG1_1;
   RS2<=READ_REG2_1;

   SHIFT: SHIFT_REG_1
      GENERIC MAP(64)
      PORT MAP (IMM_OUT1,CLK,RST,'1',IMM_OUT1_SHIFTED);

   EX_ADD: ADDER
      GENERIC MAP(64)
      PORT MAP (PC_2,IMM_OUT1_SHIFTED,'0',SUM);

   MUX_ALU: MUX_DATA
      GENERIC MAP(64)
      PORT MAP (MUX_ALU_SEL, SIGNED(IMM_OUT1), READ_DATA2_1, MUX_ALU_OUT);

   MUX_3_1: MUX_3
      GENERIC MAP(64)
      PORT MAP (FU_A, READ_DATA1_1, MUX_WB_OUT,ALU_RESULT_1_SIGNAL, READ_DATA1_2);

   MUX_3_2: MUX_3
      GENERIC MAP(64)
      PORT MAP (FU_B, MUX_ALU_OUT, MUX_WB_OUT,ALU_RESULT_1_SIGNAL, MUX_ALU_OUT_1);

  ALU_DP: ALU
      PORT MAP (READ_DATA1_2, MUX_ALU_OUT_1, ALU_OPERATION, CLK, ZERO, ALU_RESULT);

--REG EX/MEM

   REG_SUM_EX: REG
      GENERIC MAP(64)
      PORT MAP (SUM,CLK,RST,'1',SUM_1);

   REG_ALU_EX: REG_DATA
      GENERIC MAP(64)
      PORT MAP (ALU_RESULT,CLK,RST,'1',ALU_RESULT_1_SIGNAL);

   REG_READ_DATA2_EX: REG_DATA
      GENERIC MAP(64)
      PORT MAP (READ_DATA1_2,CLK,RST,'1',READ_DATA1_3);

   REG_RD_EX: REG
      GENERIC MAP(5)
      PORT MAP (RD_1,CLK,RST,'1',RD_2);  

   ALU_RESULT_1<=ALU_RESULT_1_SIGNAL;

--STAGE4

--DATA MEMORY IN TESTBENCH

--REG MEM/WB

   REG_READ_DATA_MEM: REG_DATA
      GENERIC MAP(64)
      PORT MAP (READ_DATA,CLK,RST,'1', READ_DATA_1);

   REG_ALU_MEM: REG_DATA
      GENERIC MAP(64)
      PORT MAP (ALU_RESULT_1_SIGNAL,CLK,RST,'1',ALU_RESULT_2);

   REG_RD_MEM: REG
      GENERIC MAP(5)
      PORT MAP (RD_2,CLK,RST,'1',RD_3);

--STAGE5

   MUX_WB: MUX_DATA
      GENERIC MAP(64)  
      PORT MAP (MUX_WB_SEL, READ_DATA_1, ALU_RESULT_2, MUX_WB_OUT);

END ARCHITECTURE;