LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY PC_REG IS
	PORT (
		D 				: IN UNSIGNED(63 DOWNTO 0);
		CLK,RST_N,EN 	: IN STD_LOGIC;
		Q				: OUT UNSIGNED(63 DOWNTO 0)
	);
END ENTITY;

ARCHITECTURE BEHAVIOR OF PC_REG IS

BEGIN

	PROCESS(CLK,RST_N)

	BEGIN
		IF (RST_N='0') THEN
			Q <= x"0000000000400000";
		ELSIF (CLK'EVENT AND CLK='1' AND EN='1') THEN
			Q <= D;
		END IF;

	END PROCESS;

END BEHAVIOR;