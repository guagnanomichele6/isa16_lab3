LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY FORWARDING_UNIT IS
	PORT(
		RD_2, RD_3, RS_1, RS_2: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		FU_A, FU_B: OUT STD_LOGIC_VECTOR(1 DOWNTO 0)
	);
END ENTITY;

ARCHITECTURE BEHAVIOR OF FORWARDING_UNIT IS

SIGNAL ZERO1,ZERO2,ZERO3,ZERO4: STD_LOGIC;
SIGNAL ZEROA,ZEROB: STD_LOGIC_VECTOR (1 DOWNTO 0);
COMPONENT COMPARATOR IS
	PORT(
		A, B: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		RES: OUT STD_LOGIC
	);
END COMPONENT;


BEGIN

ZERO1_1: COMPARATOR
      PORT MAP (RS_1,RD_2,ZERO1);
ZERO1_2: COMPARATOR
      PORT MAP (RS_1,RD_3,ZERO2);
ZERO2_1: COMPARATOR
      PORT MAP (RS_2,RD_2,ZERO3);
ZERO2_2: COMPARATOR
      PORT MAP (RS_2,RD_3,ZERO4);

ZEROA<=ZERO1&ZERO2;
ZEROB<=ZERO3&ZERO4;
WITH ZEROA SELECT FU_A <=
	"00" WHEN "00",
	"01" WHEN "10",
	"10" WHEN OTHERS;
WITH ZEROB SELECT FU_B <=
	"00" WHEN "00",
	"01" WHEN "10",
	"10" WHEN OTHERS;

--WITH ZERO2 SELECT FU_A(0) <=
	--'1' WHEN '1',
	--'0' WHEN OTHERS;

--WITH ZERO3 SELECT FU_B(1) <=
	--'1' WHEN '1',
	--'0' WHEN OTHERS;

--WITH ZERO4 SELECT FU_B(0) <=
	--'1' WHEN '1',
	--'0' WHEN OTHERS;


END ARCHITECTURE;