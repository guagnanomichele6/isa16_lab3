LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY ALU_CONTROL IS
	PORT(
		ALU_OP: IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		INSTR: IN STD_LOGIC_VECTOR(3 DOWNTO 0);--func(6)&func3
		ALU_OPERATION: OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END ENTITY;

ARCHITECTURE BEHAVIOR OF ALU_CONTROL IS

SIGNAL AING: STD_LOGIC_VECTOR(5 DOWNTO 0);
COMPONENT ADDER IS
        GENERIC(N:INTEGER);
	PORT (
		A 		: IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
		B 		: IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
		S 		: OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0);
		COUT 	: OUT STD_LOGIC
	);
END COMPONENT;

BEGIN

	AING<=ALU_OP&INSTR;
	WITH AING SELECT ALU_OPERATION <=
	"0010" WHEN "00-000",--ADDI
	"0000" WHEN "00-111",--ANDI
	"0011" WHEN "001101",--SRAI
	"0010" WHEN "00-010",--LW
	"0010" WHEN "01----",--U
	"0010" WHEN "100000",--ADD
	"0001" WHEN "100100", --XOR
	"0100" WHEN "100010", --SLT
	"0111" WHEN "11----", --BRANCH
	"0010" WHEN OTHERS;--ADDI?(NOP)

END ARCHITECTURE;