library verilog;
use verilog.vl_types.all;
entity tb_riscv is
end tb_riscv;
