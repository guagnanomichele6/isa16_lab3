LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY ALU IS
	PORT(
		A: IN SIGNED(63 DOWNTO 0);
		B: IN SIGNED(63 DOWNTO 0);
		ALU_OPERATION: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		CLK: IN STD_LOGIC;
		ZERO: OUT STD_LOGIC;
		ALU_RESULT: OUT SIGNED(63 DOWNTO 0)
	);
END ENTITY;

ARCHITECTURE BEHAVIOR OF ALU IS

SIGNAL ALU_RESULT_PROV_1,ALU_RESULT_PROV_2,ALU_RESULT_PROV_3,ALU_RESULT_PROV_4,ALU_RESULT_PROV_5,ZERO_SIGN: SIGNED(63 DOWNTO 0);
SIGNAL ALU_RESULT_PROV: SIGNED(63 DOWNTO 0);

COMPONENT ADD_SUB IS
        GENERIC(N:INTEGER);
	PORT (
		A 		: IN SIGNED(N-1 DOWNTO 0);
		B 		: IN SIGNED(N-1 DOWNTO 0);
		CIN		: IN STD_LOGIC;
		S 		: OUT SIGNED(N-1 DOWNTO 0)
	);
END COMPONENT;

BEGIN

ADD: ADD_SUB
      GENERIC MAP(64)
      PORT MAP (A,B,ALU_OPERATION(3),ALU_RESULT_PROV_1);

ALU_RESULT_PROV_2<=A AND B;

ALU_RESULT_PROV_3<=A XOR B;

SUB: ADD_SUB
      GENERIC MAP(64)
      PORT MAP (A,B,'1',ALU_RESULT_PROV);

    ALU_RESULT_PROV_4<=SHIFT_RIGHT(A,TO_INTEGER(UNSIGNED(B(24 DOWNTO 20))));

ALU_RESULT_PROV_5<=(63 DOWNTO 1 => '0')&ALU_RESULT_PROV(63); 

WITH ALU_OPERATION SELECT ALU_RESULT <=
	ALU_RESULT_PROV_1 WHEN "0010",--ADD
	ALU_RESULT_PROV_1 WHEN "0111",--SUB
	ALU_RESULT_PROV_2 WHEN "0000",--AND
	ALU_RESULT_PROV_3 WHEN "0001",--XOR
	ALU_RESULT_PROV_4 WHEN "0011",--SRAI
        ALU_RESULT_PROV_5 WHEN "0100",--SLT   
	ALU_RESULT_PROV_1 WHEN OTHERS;

ZERO_SIGN<= A XOR B;

WITH ZERO_SIGN SELECT ZERO <=
    '1' WHEN "0000000000000000000000000000000000000000000000000000000000000000",
    '0' WHEN OTHERS;

END ARCHITECTURE;